// see LICENSE.incore for more details on licensing terms
/*
Author: Neel Gala, neelgala@incoresemi.com
Created on: Thursday 09 April 2020 09:24:27 PM IST

*/
package apb ;

  import apb_types  :: * ;
  import apb_fabric :: * ;

  export apb_types  :: * ;
  export apb_fabric :: * ;

endpackage: apb

