// see LICENSE.incore for more details on licensing terms
/*
Author: Neel Gala, neelgala@incoresemi.com
Created on: Thursday 09 April 2020 09:52:33 PM IST

*/
package axi4 ;

  import axi4_fabric  :: * ;
  import axi4_types   :: * ;

  export axi4_fabric  :: * ;
  export axi4_types   :: * ;
endpackage: axi4

