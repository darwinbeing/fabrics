// see LICENSE.incore for more details on licensing terms
/*
Author: Neel Gala, neelgala@incoresemi.com
Created on: Thursday 09 April 2020 10:10:38 PM IST

*/
package bridges ;

  import axi2apb  :: * ;
  import axi2axil :: * ;
  import axil2apb :: * ;

  export axi2apb  :: * ;
  export axi2axil :: * ;
  export axil2apb :: * ;

endpackage: bridges

