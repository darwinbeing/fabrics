// see LICENSE.incore for more details on licensing terms
/*
Author: Babu P S, info@incoresemi.com
Created on: 25 February 2021 01:03:55 PM IST

*/
package atb ;
  import atb_types :: * ;
  import atb_components :: * ;

  export atb_types :: * ;
  export atb_components :: * ;
endpackage: atb

