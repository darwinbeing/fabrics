// see LICENSE.incore for more details on licensing terms
/*
Author: Neel Gala, neelgala@incoresemi.com
Created on: Sunday 12 April 2020 01:03:55 PM IST

*/
package axi4l ;
  import axi4l_types :: * ;
  import axi4l_fabric :: * ;

  export axi4l_types :: * ;
  export axi4l_fabric :: * ;
endpackage: axi4l

